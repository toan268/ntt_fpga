`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/22/2023 04:09:17 PM
// Design Name: 
// Module Name: NTT_GEN1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module NTT_GEN1(clk,address1,a);

	input clk;
	input [9:0] address1;
	output reg [23:0] a;
	// Declare the ROM variable
	reg [23:0] mem_ROMWRAP [895:0];


	// Initialize the ROM with $readmemb.  Put the memory contents
	// in the file dual_port_rom_init.txt.  Without this file,
	// this design will not compile.
	// See Verilog LRM 1364-2001 Section 17.2.8 for details on the
	// format of this file.

	initial 
	begin 
		mem_ROMWRAP[0] = {8'd0,8'd128,8'd1};
            mem_ROMWRAP[1] = {8'd1,8'd129,8'd1};
            mem_ROMWRAP[2] = {8'd2,8'd130,8'd1};
            mem_ROMWRAP[3] = {8'd3,8'd131,8'd1};
            mem_ROMWRAP[4] = {8'd4,8'd132,8'd1};
            mem_ROMWRAP[5] = {8'd5,8'd133,8'd1};
            mem_ROMWRAP[6] = {8'd6,8'd134,8'd1};
            mem_ROMWRAP[7] = {8'd7,8'd135,8'd1};
            mem_ROMWRAP[8] = {8'd8,8'd136,8'd1};
            mem_ROMWRAP[9] = {8'd9,8'd137,8'd1};
            mem_ROMWRAP[10] = {8'd10,8'd138,8'd1};
            mem_ROMWRAP[11] = {8'd11,8'd139,8'd1};
            mem_ROMWRAP[12] = {8'd12,8'd140,8'd1};
            mem_ROMWRAP[13] = {8'd13,8'd141,8'd1};
            mem_ROMWRAP[14] = {8'd14,8'd142,8'd1};
            mem_ROMWRAP[15] = {8'd15,8'd143,8'd1};
            mem_ROMWRAP[16] = {8'd16,8'd144,8'd1};
            mem_ROMWRAP[17] = {8'd17,8'd145,8'd1};
            mem_ROMWRAP[18] = {8'd18,8'd146,8'd1};
            mem_ROMWRAP[19] = {8'd19,8'd147,8'd1};
            mem_ROMWRAP[20] = {8'd20,8'd148,8'd1};
            mem_ROMWRAP[21] = {8'd21,8'd149,8'd1};
            mem_ROMWRAP[22] = {8'd22,8'd150,8'd1};
            mem_ROMWRAP[23] = {8'd23,8'd151,8'd1};
            mem_ROMWRAP[24] = {8'd24,8'd152,8'd1};
            mem_ROMWRAP[25] = {8'd25,8'd153,8'd1};
            mem_ROMWRAP[26] = {8'd26,8'd154,8'd1};
            mem_ROMWRAP[27] = {8'd27,8'd155,8'd1};
            mem_ROMWRAP[28] = {8'd28,8'd156,8'd1};
            mem_ROMWRAP[29] = {8'd29,8'd157,8'd1};
            mem_ROMWRAP[30] = {8'd30,8'd158,8'd1};
            mem_ROMWRAP[31] = {8'd31,8'd159,8'd1};
            mem_ROMWRAP[32] = {8'd32,8'd160,8'd1};
            mem_ROMWRAP[33] = {8'd33,8'd161,8'd1};
            mem_ROMWRAP[34] = {8'd34,8'd162,8'd1};
            mem_ROMWRAP[35] = {8'd35,8'd163,8'd1};
            mem_ROMWRAP[36] = {8'd36,8'd164,8'd1};
            mem_ROMWRAP[37] = {8'd37,8'd165,8'd1};
            mem_ROMWRAP[38] = {8'd38,8'd166,8'd1};
            mem_ROMWRAP[39] = {8'd39,8'd167,8'd1};
            mem_ROMWRAP[40] = {8'd40,8'd168,8'd1};
            mem_ROMWRAP[41] = {8'd41,8'd169,8'd1};
            mem_ROMWRAP[42] = {8'd42,8'd170,8'd1};
            mem_ROMWRAP[43] = {8'd43,8'd171,8'd1};
            mem_ROMWRAP[44] = {8'd44,8'd172,8'd1};
            mem_ROMWRAP[45] = {8'd45,8'd173,8'd1};
            mem_ROMWRAP[46] = {8'd46,8'd174,8'd1};
            mem_ROMWRAP[47] = {8'd47,8'd175,8'd1};
            mem_ROMWRAP[48] = {8'd48,8'd176,8'd1};
            mem_ROMWRAP[49] = {8'd49,8'd177,8'd1};
            mem_ROMWRAP[50] = {8'd50,8'd178,8'd1};
            mem_ROMWRAP[51] = {8'd51,8'd179,8'd1};
            mem_ROMWRAP[52] = {8'd52,8'd180,8'd1};
            mem_ROMWRAP[53] = {8'd53,8'd181,8'd1};
            mem_ROMWRAP[54] = {8'd54,8'd182,8'd1};
            mem_ROMWRAP[55] = {8'd55,8'd183,8'd1};
            mem_ROMWRAP[56] = {8'd56,8'd184,8'd1};
            mem_ROMWRAP[57] = {8'd57,8'd185,8'd1};
            mem_ROMWRAP[58] = {8'd58,8'd186,8'd1};
            mem_ROMWRAP[59] = {8'd59,8'd187,8'd1};
            mem_ROMWRAP[60] = {8'd60,8'd188,8'd1};
            mem_ROMWRAP[61] = {8'd61,8'd189,8'd1};
            mem_ROMWRAP[62] = {8'd62,8'd190,8'd1};
            mem_ROMWRAP[63] = {8'd63,8'd191,8'd1};
            mem_ROMWRAP[64] = {8'd64,8'd192,8'd1};
            mem_ROMWRAP[65] = {8'd65,8'd193,8'd1};
            mem_ROMWRAP[66] = {8'd66,8'd194,8'd1};
            mem_ROMWRAP[67] = {8'd67,8'd195,8'd1};
            mem_ROMWRAP[68] = {8'd68,8'd196,8'd1};
            mem_ROMWRAP[69] = {8'd69,8'd197,8'd1};
            mem_ROMWRAP[70] = {8'd70,8'd198,8'd1};
            mem_ROMWRAP[71] = {8'd71,8'd199,8'd1};
            mem_ROMWRAP[72] = {8'd72,8'd200,8'd1};
            mem_ROMWRAP[73] = {8'd73,8'd201,8'd1};
            mem_ROMWRAP[74] = {8'd74,8'd202,8'd1};
            mem_ROMWRAP[75] = {8'd75,8'd203,8'd1};
            mem_ROMWRAP[76] = {8'd76,8'd204,8'd1};
            mem_ROMWRAP[77] = {8'd77,8'd205,8'd1};
            mem_ROMWRAP[78] = {8'd78,8'd206,8'd1};
            mem_ROMWRAP[79] = {8'd79,8'd207,8'd1};
            mem_ROMWRAP[80] = {8'd80,8'd208,8'd1};
            mem_ROMWRAP[81] = {8'd81,8'd209,8'd1};
            mem_ROMWRAP[82] = {8'd82,8'd210,8'd1};
            mem_ROMWRAP[83] = {8'd83,8'd211,8'd1};
            mem_ROMWRAP[84] = {8'd84,8'd212,8'd1};
            mem_ROMWRAP[85] = {8'd85,8'd213,8'd1};
            mem_ROMWRAP[86] = {8'd86,8'd214,8'd1};
            mem_ROMWRAP[87] = {8'd87,8'd215,8'd1};
            mem_ROMWRAP[88] = {8'd88,8'd216,8'd1};
            mem_ROMWRAP[89] = {8'd89,8'd217,8'd1};
            mem_ROMWRAP[90] = {8'd90,8'd218,8'd1};
            mem_ROMWRAP[91] = {8'd91,8'd219,8'd1};
            mem_ROMWRAP[92] = {8'd92,8'd220,8'd1};
            mem_ROMWRAP[93] = {8'd93,8'd221,8'd1};
            mem_ROMWRAP[94] = {8'd94,8'd222,8'd1};
            mem_ROMWRAP[95] = {8'd95,8'd223,8'd1};
            mem_ROMWRAP[96] = {8'd96,8'd224,8'd1};
            mem_ROMWRAP[97] = {8'd97,8'd225,8'd1};
            mem_ROMWRAP[98] = {8'd98,8'd226,8'd1};
            mem_ROMWRAP[99] = {8'd99,8'd227,8'd1};
            mem_ROMWRAP[100] = {8'd100,8'd228,8'd1};
            mem_ROMWRAP[101] = {8'd101,8'd229,8'd1};
            mem_ROMWRAP[102] = {8'd102,8'd230,8'd1};
            mem_ROMWRAP[103] = {8'd103,8'd231,8'd1};
            mem_ROMWRAP[104] = {8'd104,8'd232,8'd1};
            mem_ROMWRAP[105] = {8'd105,8'd233,8'd1};
            mem_ROMWRAP[106] = {8'd106,8'd234,8'd1};
            mem_ROMWRAP[107] = {8'd107,8'd235,8'd1};
            mem_ROMWRAP[108] = {8'd108,8'd236,8'd1};
            mem_ROMWRAP[109] = {8'd109,8'd237,8'd1};
            mem_ROMWRAP[110] = {8'd110,8'd238,8'd1};
            mem_ROMWRAP[111] = {8'd111,8'd239,8'd1};
            mem_ROMWRAP[112] = {8'd112,8'd240,8'd1};
            mem_ROMWRAP[113] = {8'd113,8'd241,8'd1};
            mem_ROMWRAP[114] = {8'd114,8'd242,8'd1};
            mem_ROMWRAP[115] = {8'd115,8'd243,8'd1};
            mem_ROMWRAP[116] = {8'd116,8'd244,8'd1};
            mem_ROMWRAP[117] = {8'd117,8'd245,8'd1};
            mem_ROMWRAP[118] = {8'd118,8'd246,8'd1};
            mem_ROMWRAP[119] = {8'd119,8'd247,8'd1};
            mem_ROMWRAP[120] = {8'd120,8'd248,8'd1};
            mem_ROMWRAP[121] = {8'd121,8'd249,8'd1};
            mem_ROMWRAP[122] = {8'd122,8'd250,8'd1};
            mem_ROMWRAP[123] = {8'd123,8'd251,8'd1};
            mem_ROMWRAP[124] = {8'd124,8'd252,8'd1};
            mem_ROMWRAP[125] = {8'd125,8'd253,8'd1};
            mem_ROMWRAP[126] = {8'd126,8'd254,8'd1};
            mem_ROMWRAP[127] = {8'd127,8'd255,8'd1};
            mem_ROMWRAP[128] = {8'd0,8'd64,8'd2};
            mem_ROMWRAP[129] = {8'd1,8'd65,8'd2};
            mem_ROMWRAP[130] = {8'd2,8'd66,8'd2};
            mem_ROMWRAP[131] = {8'd3,8'd67,8'd2};
            mem_ROMWRAP[132] = {8'd4,8'd68,8'd2};
            mem_ROMWRAP[133] = {8'd5,8'd69,8'd2};
            mem_ROMWRAP[134] = {8'd6,8'd70,8'd2};
            mem_ROMWRAP[135] = {8'd7,8'd71,8'd2};
            mem_ROMWRAP[136] = {8'd8,8'd72,8'd2};
            mem_ROMWRAP[137] = {8'd9,8'd73,8'd2};
            mem_ROMWRAP[138] = {8'd10,8'd74,8'd2};
            mem_ROMWRAP[139] = {8'd11,8'd75,8'd2};
            mem_ROMWRAP[140] = {8'd12,8'd76,8'd2};
            mem_ROMWRAP[141] = {8'd13,8'd77,8'd2};
            mem_ROMWRAP[142] = {8'd14,8'd78,8'd2};
            mem_ROMWRAP[143] = {8'd15,8'd79,8'd2};
            mem_ROMWRAP[144] = {8'd16,8'd80,8'd2};
            mem_ROMWRAP[145] = {8'd17,8'd81,8'd2};
            mem_ROMWRAP[146] = {8'd18,8'd82,8'd2};
            mem_ROMWRAP[147] = {8'd19,8'd83,8'd2};
            mem_ROMWRAP[148] = {8'd20,8'd84,8'd2};
            mem_ROMWRAP[149] = {8'd21,8'd85,8'd2};
            mem_ROMWRAP[150] = {8'd22,8'd86,8'd2};
            mem_ROMWRAP[151] = {8'd23,8'd87,8'd2};
            mem_ROMWRAP[152] = {8'd24,8'd88,8'd2};
            mem_ROMWRAP[153] = {8'd25,8'd89,8'd2};
            mem_ROMWRAP[154] = {8'd26,8'd90,8'd2};
            mem_ROMWRAP[155] = {8'd27,8'd91,8'd2};
            mem_ROMWRAP[156] = {8'd28,8'd92,8'd2};
            mem_ROMWRAP[157] = {8'd29,8'd93,8'd2};
            mem_ROMWRAP[158] = {8'd30,8'd94,8'd2};
            mem_ROMWRAP[159] = {8'd31,8'd95,8'd2};
            mem_ROMWRAP[160] = {8'd32,8'd96,8'd2};
            mem_ROMWRAP[161] = {8'd33,8'd97,8'd2};
            mem_ROMWRAP[162] = {8'd34,8'd98,8'd2};
            mem_ROMWRAP[163] = {8'd35,8'd99,8'd2};
            mem_ROMWRAP[164] = {8'd36,8'd100,8'd2};
            mem_ROMWRAP[165] = {8'd37,8'd101,8'd2};
            mem_ROMWRAP[166] = {8'd38,8'd102,8'd2};
            mem_ROMWRAP[167] = {8'd39,8'd103,8'd2};
            mem_ROMWRAP[168] = {8'd40,8'd104,8'd2};
            mem_ROMWRAP[169] = {8'd41,8'd105,8'd2};
            mem_ROMWRAP[170] = {8'd42,8'd106,8'd2};
            mem_ROMWRAP[171] = {8'd43,8'd107,8'd2};
            mem_ROMWRAP[172] = {8'd44,8'd108,8'd2};
            mem_ROMWRAP[173] = {8'd45,8'd109,8'd2};
            mem_ROMWRAP[174] = {8'd46,8'd110,8'd2};
            mem_ROMWRAP[175] = {8'd47,8'd111,8'd2};
            mem_ROMWRAP[176] = {8'd48,8'd112,8'd2};
            mem_ROMWRAP[177] = {8'd49,8'd113,8'd2};
            mem_ROMWRAP[178] = {8'd50,8'd114,8'd2};
            mem_ROMWRAP[179] = {8'd51,8'd115,8'd2};
            mem_ROMWRAP[180] = {8'd52,8'd116,8'd2};
            mem_ROMWRAP[181] = {8'd53,8'd117,8'd2};
            mem_ROMWRAP[182] = {8'd54,8'd118,8'd2};
            mem_ROMWRAP[183] = {8'd55,8'd119,8'd2};
            mem_ROMWRAP[184] = {8'd56,8'd120,8'd2};
            mem_ROMWRAP[185] = {8'd57,8'd121,8'd2};
            mem_ROMWRAP[186] = {8'd58,8'd122,8'd2};
            mem_ROMWRAP[187] = {8'd59,8'd123,8'd2};
            mem_ROMWRAP[188] = {8'd60,8'd124,8'd2};
            mem_ROMWRAP[189] = {8'd61,8'd125,8'd2};
            mem_ROMWRAP[190] = {8'd62,8'd126,8'd2};
            mem_ROMWRAP[191] = {8'd63,8'd127,8'd2};
            mem_ROMWRAP[192] = {8'd128,8'd192,8'd3};
            mem_ROMWRAP[193] = {8'd129,8'd193,8'd3};
            mem_ROMWRAP[194] = {8'd130,8'd194,8'd3};
            mem_ROMWRAP[195] = {8'd131,8'd195,8'd3};
            mem_ROMWRAP[196] = {8'd132,8'd196,8'd3};
            mem_ROMWRAP[197] = {8'd133,8'd197,8'd3};
            mem_ROMWRAP[198] = {8'd134,8'd198,8'd3};
            mem_ROMWRAP[199] = {8'd135,8'd199,8'd3};
            mem_ROMWRAP[200] = {8'd136,8'd200,8'd3};
            mem_ROMWRAP[201] = {8'd137,8'd201,8'd3};
            mem_ROMWRAP[202] = {8'd138,8'd202,8'd3};
            mem_ROMWRAP[203] = {8'd139,8'd203,8'd3};
            mem_ROMWRAP[204] = {8'd140,8'd204,8'd3};
            mem_ROMWRAP[205] = {8'd141,8'd205,8'd3};
            mem_ROMWRAP[206] = {8'd142,8'd206,8'd3};
            mem_ROMWRAP[207] = {8'd143,8'd207,8'd3};
            mem_ROMWRAP[208] = {8'd144,8'd208,8'd3};
            mem_ROMWRAP[209] = {8'd145,8'd209,8'd3};
            mem_ROMWRAP[210] = {8'd146,8'd210,8'd3};
            mem_ROMWRAP[211] = {8'd147,8'd211,8'd3};
            mem_ROMWRAP[212] = {8'd148,8'd212,8'd3};
            mem_ROMWRAP[213] = {8'd149,8'd213,8'd3};
            mem_ROMWRAP[214] = {8'd150,8'd214,8'd3};
            mem_ROMWRAP[215] = {8'd151,8'd215,8'd3};
            mem_ROMWRAP[216] = {8'd152,8'd216,8'd3};
            mem_ROMWRAP[217] = {8'd153,8'd217,8'd3};
            mem_ROMWRAP[218] = {8'd154,8'd218,8'd3};
            mem_ROMWRAP[219] = {8'd155,8'd219,8'd3};
            mem_ROMWRAP[220] = {8'd156,8'd220,8'd3};
            mem_ROMWRAP[221] = {8'd157,8'd221,8'd3};
            mem_ROMWRAP[222] = {8'd158,8'd222,8'd3};
            mem_ROMWRAP[223] = {8'd159,8'd223,8'd3};
            mem_ROMWRAP[224] = {8'd160,8'd224,8'd3};
            mem_ROMWRAP[225] = {8'd161,8'd225,8'd3};
            mem_ROMWRAP[226] = {8'd162,8'd226,8'd3};
            mem_ROMWRAP[227] = {8'd163,8'd227,8'd3};
            mem_ROMWRAP[228] = {8'd164,8'd228,8'd3};
            mem_ROMWRAP[229] = {8'd165,8'd229,8'd3};
            mem_ROMWRAP[230] = {8'd166,8'd230,8'd3};
            mem_ROMWRAP[231] = {8'd167,8'd231,8'd3};
            mem_ROMWRAP[232] = {8'd168,8'd232,8'd3};
            mem_ROMWRAP[233] = {8'd169,8'd233,8'd3};
            mem_ROMWRAP[234] = {8'd170,8'd234,8'd3};
            mem_ROMWRAP[235] = {8'd171,8'd235,8'd3};
            mem_ROMWRAP[236] = {8'd172,8'd236,8'd3};
            mem_ROMWRAP[237] = {8'd173,8'd237,8'd3};
            mem_ROMWRAP[238] = {8'd174,8'd238,8'd3};
            mem_ROMWRAP[239] = {8'd175,8'd239,8'd3};
            mem_ROMWRAP[240] = {8'd176,8'd240,8'd3};
            mem_ROMWRAP[241] = {8'd177,8'd241,8'd3};
            mem_ROMWRAP[242] = {8'd178,8'd242,8'd3};
            mem_ROMWRAP[243] = {8'd179,8'd243,8'd3};
            mem_ROMWRAP[244] = {8'd180,8'd244,8'd3};
            mem_ROMWRAP[245] = {8'd181,8'd245,8'd3};
            mem_ROMWRAP[246] = {8'd182,8'd246,8'd3};
            mem_ROMWRAP[247] = {8'd183,8'd247,8'd3};
            mem_ROMWRAP[248] = {8'd184,8'd248,8'd3};
            mem_ROMWRAP[249] = {8'd185,8'd249,8'd3};
            mem_ROMWRAP[250] = {8'd186,8'd250,8'd3};
            mem_ROMWRAP[251] = {8'd187,8'd251,8'd3};
            mem_ROMWRAP[252] = {8'd188,8'd252,8'd3};
            mem_ROMWRAP[253] = {8'd189,8'd253,8'd3};
            mem_ROMWRAP[254] = {8'd190,8'd254,8'd3};
            mem_ROMWRAP[255] = {8'd191,8'd255,8'd3};
            mem_ROMWRAP[256] = {8'd0,8'd32,8'd4};
            mem_ROMWRAP[257] = {8'd1,8'd33,8'd4};
            mem_ROMWRAP[258] = {8'd2,8'd34,8'd4};
            mem_ROMWRAP[259] = {8'd3,8'd35,8'd4};
            mem_ROMWRAP[260] = {8'd4,8'd36,8'd4};
            mem_ROMWRAP[261] = {8'd5,8'd37,8'd4};
            mem_ROMWRAP[262] = {8'd6,8'd38,8'd4};
            mem_ROMWRAP[263] = {8'd7,8'd39,8'd4};
            mem_ROMWRAP[264] = {8'd8,8'd40,8'd4};
            mem_ROMWRAP[265] = {8'd9,8'd41,8'd4};
            mem_ROMWRAP[266] = {8'd10,8'd42,8'd4};
            mem_ROMWRAP[267] = {8'd11,8'd43,8'd4};
            mem_ROMWRAP[268] = {8'd12,8'd44,8'd4};
            mem_ROMWRAP[269] = {8'd13,8'd45,8'd4};
            mem_ROMWRAP[270] = {8'd14,8'd46,8'd4};
            mem_ROMWRAP[271] = {8'd15,8'd47,8'd4};
            mem_ROMWRAP[272] = {8'd16,8'd48,8'd4};
            mem_ROMWRAP[273] = {8'd17,8'd49,8'd4};
            mem_ROMWRAP[274] = {8'd18,8'd50,8'd4};
            mem_ROMWRAP[275] = {8'd19,8'd51,8'd4};
            mem_ROMWRAP[276] = {8'd20,8'd52,8'd4};
            mem_ROMWRAP[277] = {8'd21,8'd53,8'd4};
            mem_ROMWRAP[278] = {8'd22,8'd54,8'd4};
            mem_ROMWRAP[279] = {8'd23,8'd55,8'd4};
            mem_ROMWRAP[280] = {8'd24,8'd56,8'd4};
            mem_ROMWRAP[281] = {8'd25,8'd57,8'd4};
            mem_ROMWRAP[282] = {8'd26,8'd58,8'd4};
            mem_ROMWRAP[283] = {8'd27,8'd59,8'd4};
            mem_ROMWRAP[284] = {8'd28,8'd60,8'd4};
            mem_ROMWRAP[285] = {8'd29,8'd61,8'd4};
            mem_ROMWRAP[286] = {8'd30,8'd62,8'd4};
            mem_ROMWRAP[287] = {8'd31,8'd63,8'd4};
            mem_ROMWRAP[288] = {8'd64,8'd96,8'd5};
            mem_ROMWRAP[289] = {8'd65,8'd97,8'd5};
            mem_ROMWRAP[290] = {8'd66,8'd98,8'd5};
            mem_ROMWRAP[291] = {8'd67,8'd99,8'd5};
            mem_ROMWRAP[292] = {8'd68,8'd100,8'd5};
            mem_ROMWRAP[293] = {8'd69,8'd101,8'd5};
            mem_ROMWRAP[294] = {8'd70,8'd102,8'd5};
            mem_ROMWRAP[295] = {8'd71,8'd103,8'd5};
            mem_ROMWRAP[296] = {8'd72,8'd104,8'd5};
            mem_ROMWRAP[297] = {8'd73,8'd105,8'd5};
            mem_ROMWRAP[298] = {8'd74,8'd106,8'd5};
            mem_ROMWRAP[299] = {8'd75,8'd107,8'd5};
            mem_ROMWRAP[300] = {8'd76,8'd108,8'd5};
            mem_ROMWRAP[301] = {8'd77,8'd109,8'd5};
            mem_ROMWRAP[302] = {8'd78,8'd110,8'd5};
            mem_ROMWRAP[303] = {8'd79,8'd111,8'd5};
            mem_ROMWRAP[304] = {8'd80,8'd112,8'd5};
            mem_ROMWRAP[305] = {8'd81,8'd113,8'd5};
            mem_ROMWRAP[306] = {8'd82,8'd114,8'd5};
            mem_ROMWRAP[307] = {8'd83,8'd115,8'd5};
            mem_ROMWRAP[308] = {8'd84,8'd116,8'd5};
            mem_ROMWRAP[309] = {8'd85,8'd117,8'd5};
            mem_ROMWRAP[310] = {8'd86,8'd118,8'd5};
            mem_ROMWRAP[311] = {8'd87,8'd119,8'd5};
            mem_ROMWRAP[312] = {8'd88,8'd120,8'd5};
            mem_ROMWRAP[313] = {8'd89,8'd121,8'd5};
            mem_ROMWRAP[314] = {8'd90,8'd122,8'd5};
            mem_ROMWRAP[315] = {8'd91,8'd123,8'd5};
            mem_ROMWRAP[316] = {8'd92,8'd124,8'd5};
            mem_ROMWRAP[317] = {8'd93,8'd125,8'd5};
            mem_ROMWRAP[318] = {8'd94,8'd126,8'd5};
            mem_ROMWRAP[319] = {8'd95,8'd127,8'd5};
            mem_ROMWRAP[320] = {8'd128,8'd160,8'd6};
            mem_ROMWRAP[321] = {8'd129,8'd161,8'd6};
            mem_ROMWRAP[322] = {8'd130,8'd162,8'd6};
            mem_ROMWRAP[323] = {8'd131,8'd163,8'd6};
            mem_ROMWRAP[324] = {8'd132,8'd164,8'd6};
            mem_ROMWRAP[325] = {8'd133,8'd165,8'd6};
            mem_ROMWRAP[326] = {8'd134,8'd166,8'd6};
            mem_ROMWRAP[327] = {8'd135,8'd167,8'd6};
            mem_ROMWRAP[328] = {8'd136,8'd168,8'd6};
            mem_ROMWRAP[329] = {8'd137,8'd169,8'd6};
            mem_ROMWRAP[330] = {8'd138,8'd170,8'd6};
            mem_ROMWRAP[331] = {8'd139,8'd171,8'd6};
            mem_ROMWRAP[332] = {8'd140,8'd172,8'd6};
            mem_ROMWRAP[333] = {8'd141,8'd173,8'd6};
            mem_ROMWRAP[334] = {8'd142,8'd174,8'd6};
            mem_ROMWRAP[335] = {8'd143,8'd175,8'd6};
            mem_ROMWRAP[336] = {8'd144,8'd176,8'd6};
            mem_ROMWRAP[337] = {8'd145,8'd177,8'd6};
            mem_ROMWRAP[338] = {8'd146,8'd178,8'd6};
            mem_ROMWRAP[339] = {8'd147,8'd179,8'd6};
            mem_ROMWRAP[340] = {8'd148,8'd180,8'd6};
            mem_ROMWRAP[341] = {8'd149,8'd181,8'd6};
            mem_ROMWRAP[342] = {8'd150,8'd182,8'd6};
            mem_ROMWRAP[343] = {8'd151,8'd183,8'd6};
            mem_ROMWRAP[344] = {8'd152,8'd184,8'd6};
            mem_ROMWRAP[345] = {8'd153,8'd185,8'd6};
            mem_ROMWRAP[346] = {8'd154,8'd186,8'd6};
            mem_ROMWRAP[347] = {8'd155,8'd187,8'd6};
            mem_ROMWRAP[348] = {8'd156,8'd188,8'd6};
            mem_ROMWRAP[349] = {8'd157,8'd189,8'd6};
            mem_ROMWRAP[350] = {8'd158,8'd190,8'd6};
            mem_ROMWRAP[351] = {8'd159,8'd191,8'd6};
            mem_ROMWRAP[352] = {8'd192,8'd224,8'd7};
            mem_ROMWRAP[353] = {8'd193,8'd225,8'd7};
            mem_ROMWRAP[354] = {8'd194,8'd226,8'd7};
            mem_ROMWRAP[355] = {8'd195,8'd227,8'd7};
            mem_ROMWRAP[356] = {8'd196,8'd228,8'd7};
            mem_ROMWRAP[357] = {8'd197,8'd229,8'd7};
            mem_ROMWRAP[358] = {8'd198,8'd230,8'd7};
            mem_ROMWRAP[359] = {8'd199,8'd231,8'd7};
            mem_ROMWRAP[360] = {8'd200,8'd232,8'd7};
            mem_ROMWRAP[361] = {8'd201,8'd233,8'd7};
            mem_ROMWRAP[362] = {8'd202,8'd234,8'd7};
            mem_ROMWRAP[363] = {8'd203,8'd235,8'd7};
            mem_ROMWRAP[364] = {8'd204,8'd236,8'd7};
            mem_ROMWRAP[365] = {8'd205,8'd237,8'd7};
            mem_ROMWRAP[366] = {8'd206,8'd238,8'd7};
            mem_ROMWRAP[367] = {8'd207,8'd239,8'd7};
            mem_ROMWRAP[368] = {8'd208,8'd240,8'd7};
            mem_ROMWRAP[369] = {8'd209,8'd241,8'd7};
            mem_ROMWRAP[370] = {8'd210,8'd242,8'd7};
            mem_ROMWRAP[371] = {8'd211,8'd243,8'd7};
            mem_ROMWRAP[372] = {8'd212,8'd244,8'd7};
            mem_ROMWRAP[373] = {8'd213,8'd245,8'd7};
            mem_ROMWRAP[374] = {8'd214,8'd246,8'd7};
            mem_ROMWRAP[375] = {8'd215,8'd247,8'd7};
            mem_ROMWRAP[376] = {8'd216,8'd248,8'd7};
            mem_ROMWRAP[377] = {8'd217,8'd249,8'd7};
            mem_ROMWRAP[378] = {8'd218,8'd250,8'd7};
            mem_ROMWRAP[379] = {8'd219,8'd251,8'd7};
            mem_ROMWRAP[380] = {8'd220,8'd252,8'd7};
            mem_ROMWRAP[381] = {8'd221,8'd253,8'd7};
            mem_ROMWRAP[382] = {8'd222,8'd254,8'd7};
            mem_ROMWRAP[383] = {8'd223,8'd255,8'd7};
            mem_ROMWRAP[384] = {8'd0,8'd16,8'd8};
            mem_ROMWRAP[385] = {8'd1,8'd17,8'd8};
            mem_ROMWRAP[386] = {8'd2,8'd18,8'd8};
            mem_ROMWRAP[387] = {8'd3,8'd19,8'd8};
            mem_ROMWRAP[388] = {8'd4,8'd20,8'd8};
            mem_ROMWRAP[389] = {8'd5,8'd21,8'd8};
            mem_ROMWRAP[390] = {8'd6,8'd22,8'd8};
            mem_ROMWRAP[391] = {8'd7,8'd23,8'd8};
            mem_ROMWRAP[392] = {8'd8,8'd24,8'd8};
            mem_ROMWRAP[393] = {8'd9,8'd25,8'd8};
            mem_ROMWRAP[394] = {8'd10,8'd26,8'd8};
            mem_ROMWRAP[395] = {8'd11,8'd27,8'd8};
            mem_ROMWRAP[396] = {8'd12,8'd28,8'd8};
            mem_ROMWRAP[397] = {8'd13,8'd29,8'd8};
            mem_ROMWRAP[398] = {8'd14,8'd30,8'd8};
            mem_ROMWRAP[399] = {8'd15,8'd31,8'd8};
            mem_ROMWRAP[400] = {8'd32,8'd48,8'd9};
            mem_ROMWRAP[401] = {8'd33,8'd49,8'd9};
            mem_ROMWRAP[402] = {8'd34,8'd50,8'd9};
            mem_ROMWRAP[403] = {8'd35,8'd51,8'd9};
            mem_ROMWRAP[404] = {8'd36,8'd52,8'd9};
            mem_ROMWRAP[405] = {8'd37,8'd53,8'd9};
            mem_ROMWRAP[406] = {8'd38,8'd54,8'd9};
            mem_ROMWRAP[407] = {8'd39,8'd55,8'd9};
            mem_ROMWRAP[408] = {8'd40,8'd56,8'd9};
            mem_ROMWRAP[409] = {8'd41,8'd57,8'd9};
            mem_ROMWRAP[410] = {8'd42,8'd58,8'd9};
            mem_ROMWRAP[411] = {8'd43,8'd59,8'd9};
            mem_ROMWRAP[412] = {8'd44,8'd60,8'd9};
            mem_ROMWRAP[413] = {8'd45,8'd61,8'd9};
            mem_ROMWRAP[414] = {8'd46,8'd62,8'd9};
            mem_ROMWRAP[415] = {8'd47,8'd63,8'd9};
            mem_ROMWRAP[416] = {8'd64,8'd80,8'd10};
            mem_ROMWRAP[417] = {8'd65,8'd81,8'd10};
            mem_ROMWRAP[418] = {8'd66,8'd82,8'd10};
            mem_ROMWRAP[419] = {8'd67,8'd83,8'd10};
            mem_ROMWRAP[420] = {8'd68,8'd84,8'd10};
            mem_ROMWRAP[421] = {8'd69,8'd85,8'd10};
            mem_ROMWRAP[422] = {8'd70,8'd86,8'd10};
            mem_ROMWRAP[423] = {8'd71,8'd87,8'd10};
            mem_ROMWRAP[424] = {8'd72,8'd88,8'd10};
            mem_ROMWRAP[425] = {8'd73,8'd89,8'd10};
            mem_ROMWRAP[426] = {8'd74,8'd90,8'd10};
            mem_ROMWRAP[427] = {8'd75,8'd91,8'd10};
            mem_ROMWRAP[428] = {8'd76,8'd92,8'd10};
            mem_ROMWRAP[429] = {8'd77,8'd93,8'd10};
            mem_ROMWRAP[430] = {8'd78,8'd94,8'd10};
            mem_ROMWRAP[431] = {8'd79,8'd95,8'd10};
            mem_ROMWRAP[432] = {8'd96,8'd112,8'd11};
            mem_ROMWRAP[433] = {8'd97,8'd113,8'd11};
            mem_ROMWRAP[434] = {8'd98,8'd114,8'd11};
            mem_ROMWRAP[435] = {8'd99,8'd115,8'd11};
            mem_ROMWRAP[436] = {8'd100,8'd116,8'd11};
            mem_ROMWRAP[437] = {8'd101,8'd117,8'd11};
            mem_ROMWRAP[438] = {8'd102,8'd118,8'd11};
            mem_ROMWRAP[439] = {8'd103,8'd119,8'd11};
            mem_ROMWRAP[440] = {8'd104,8'd120,8'd11};
            mem_ROMWRAP[441] = {8'd105,8'd121,8'd11};
            mem_ROMWRAP[442] = {8'd106,8'd122,8'd11};
            mem_ROMWRAP[443] = {8'd107,8'd123,8'd11};
            mem_ROMWRAP[444] = {8'd108,8'd124,8'd11};
            mem_ROMWRAP[445] = {8'd109,8'd125,8'd11};
            mem_ROMWRAP[446] = {8'd110,8'd126,8'd11};
            mem_ROMWRAP[447] = {8'd111,8'd127,8'd11};
            mem_ROMWRAP[448] = {8'd128,8'd144,8'd12};
            mem_ROMWRAP[449] = {8'd129,8'd145,8'd12};
            mem_ROMWRAP[450] = {8'd130,8'd146,8'd12};
            mem_ROMWRAP[451] = {8'd131,8'd147,8'd12};
            mem_ROMWRAP[452] = {8'd132,8'd148,8'd12};
            mem_ROMWRAP[453] = {8'd133,8'd149,8'd12};
            mem_ROMWRAP[454] = {8'd134,8'd150,8'd12};
            mem_ROMWRAP[455] = {8'd135,8'd151,8'd12};
            mem_ROMWRAP[456] = {8'd136,8'd152,8'd12};
            mem_ROMWRAP[457] = {8'd137,8'd153,8'd12};
            mem_ROMWRAP[458] = {8'd138,8'd154,8'd12};
            mem_ROMWRAP[459] = {8'd139,8'd155,8'd12};
            mem_ROMWRAP[460] = {8'd140,8'd156,8'd12};
            mem_ROMWRAP[461] = {8'd141,8'd157,8'd12};
            mem_ROMWRAP[462] = {8'd142,8'd158,8'd12};
            mem_ROMWRAP[463] = {8'd143,8'd159,8'd12};
            mem_ROMWRAP[464] = {8'd160,8'd176,8'd13};
            mem_ROMWRAP[465] = {8'd161,8'd177,8'd13};
            mem_ROMWRAP[466] = {8'd162,8'd178,8'd13};
            mem_ROMWRAP[467] = {8'd163,8'd179,8'd13};
            mem_ROMWRAP[468] = {8'd164,8'd180,8'd13};
            mem_ROMWRAP[469] = {8'd165,8'd181,8'd13};
            mem_ROMWRAP[470] = {8'd166,8'd182,8'd13};
            mem_ROMWRAP[471] = {8'd167,8'd183,8'd13};
            mem_ROMWRAP[472] = {8'd168,8'd184,8'd13};
            mem_ROMWRAP[473] = {8'd169,8'd185,8'd13};
            mem_ROMWRAP[474] = {8'd170,8'd186,8'd13};
            mem_ROMWRAP[475] = {8'd171,8'd187,8'd13};
            mem_ROMWRAP[476] = {8'd172,8'd188,8'd13};
            mem_ROMWRAP[477] = {8'd173,8'd189,8'd13};
            mem_ROMWRAP[478] = {8'd174,8'd190,8'd13};
            mem_ROMWRAP[479] = {8'd175,8'd191,8'd13};
            mem_ROMWRAP[480] = {8'd192,8'd208,8'd14};
            mem_ROMWRAP[481] = {8'd193,8'd209,8'd14};
            mem_ROMWRAP[482] = {8'd194,8'd210,8'd14};
            mem_ROMWRAP[483] = {8'd195,8'd211,8'd14};
            mem_ROMWRAP[484] = {8'd196,8'd212,8'd14};
            mem_ROMWRAP[485] = {8'd197,8'd213,8'd14};
            mem_ROMWRAP[486] = {8'd198,8'd214,8'd14};
            mem_ROMWRAP[487] = {8'd199,8'd215,8'd14};
            mem_ROMWRAP[488] = {8'd200,8'd216,8'd14};
            mem_ROMWRAP[489] = {8'd201,8'd217,8'd14};
            mem_ROMWRAP[490] = {8'd202,8'd218,8'd14};
            mem_ROMWRAP[491] = {8'd203,8'd219,8'd14};
            mem_ROMWRAP[492] = {8'd204,8'd220,8'd14};
            mem_ROMWRAP[493] = {8'd205,8'd221,8'd14};
            mem_ROMWRAP[494] = {8'd206,8'd222,8'd14};
            mem_ROMWRAP[495] = {8'd207,8'd223,8'd14};
            mem_ROMWRAP[496] = {8'd224,8'd240,8'd15};
            mem_ROMWRAP[497] = {8'd225,8'd241,8'd15};
            mem_ROMWRAP[498] = {8'd226,8'd242,8'd15};
            mem_ROMWRAP[499] = {8'd227,8'd243,8'd15};
            mem_ROMWRAP[500] = {8'd228,8'd244,8'd15};
            mem_ROMWRAP[501] = {8'd229,8'd245,8'd15};
            mem_ROMWRAP[502] = {8'd230,8'd246,8'd15};
            mem_ROMWRAP[503] = {8'd231,8'd247,8'd15};
            mem_ROMWRAP[504] = {8'd232,8'd248,8'd15};
            mem_ROMWRAP[505] = {8'd233,8'd249,8'd15};
            mem_ROMWRAP[506] = {8'd234,8'd250,8'd15};
            mem_ROMWRAP[507] = {8'd235,8'd251,8'd15};
            mem_ROMWRAP[508] = {8'd236,8'd252,8'd15};
            mem_ROMWRAP[509] = {8'd237,8'd253,8'd15};
            mem_ROMWRAP[510] = {8'd238,8'd254,8'd15};
            mem_ROMWRAP[511] = {8'd239,8'd255,8'd15};
            mem_ROMWRAP[512] = {8'd0,8'd8,8'd16};
            mem_ROMWRAP[513] = {8'd1,8'd9,8'd16};
            mem_ROMWRAP[514] = {8'd2,8'd10,8'd16};
            mem_ROMWRAP[515] = {8'd3,8'd11,8'd16};
            mem_ROMWRAP[516] = {8'd4,8'd12,8'd16};
            mem_ROMWRAP[517] = {8'd5,8'd13,8'd16};
            mem_ROMWRAP[518] = {8'd6,8'd14,8'd16};
            mem_ROMWRAP[519] = {8'd7,8'd15,8'd16};
            mem_ROMWRAP[520] = {8'd16,8'd24,8'd17};
            mem_ROMWRAP[521] = {8'd17,8'd25,8'd17};
            mem_ROMWRAP[522] = {8'd18,8'd26,8'd17};
            mem_ROMWRAP[523] = {8'd19,8'd27,8'd17};
            mem_ROMWRAP[524] = {8'd20,8'd28,8'd17};
            mem_ROMWRAP[525] = {8'd21,8'd29,8'd17};
            mem_ROMWRAP[526] = {8'd22,8'd30,8'd17};
            mem_ROMWRAP[527] = {8'd23,8'd31,8'd17};
            mem_ROMWRAP[528] = {8'd32,8'd40,8'd18};
            mem_ROMWRAP[529] = {8'd33,8'd41,8'd18};
            mem_ROMWRAP[530] = {8'd34,8'd42,8'd18};
            mem_ROMWRAP[531] = {8'd35,8'd43,8'd18};
            mem_ROMWRAP[532] = {8'd36,8'd44,8'd18};
            mem_ROMWRAP[533] = {8'd37,8'd45,8'd18};
            mem_ROMWRAP[534] = {8'd38,8'd46,8'd18};
            mem_ROMWRAP[535] = {8'd39,8'd47,8'd18};
            mem_ROMWRAP[536] = {8'd48,8'd56,8'd19};
            mem_ROMWRAP[537] = {8'd49,8'd57,8'd19};
            mem_ROMWRAP[538] = {8'd50,8'd58,8'd19};
            mem_ROMWRAP[539] = {8'd51,8'd59,8'd19};
            mem_ROMWRAP[540] = {8'd52,8'd60,8'd19};
            mem_ROMWRAP[541] = {8'd53,8'd61,8'd19};
            mem_ROMWRAP[542] = {8'd54,8'd62,8'd19};
            mem_ROMWRAP[543] = {8'd55,8'd63,8'd19};
            mem_ROMWRAP[544] = {8'd64,8'd72,8'd20};
            mem_ROMWRAP[545] = {8'd65,8'd73,8'd20};
            mem_ROMWRAP[546] = {8'd66,8'd74,8'd20};
            mem_ROMWRAP[547] = {8'd67,8'd75,8'd20};
            mem_ROMWRAP[548] = {8'd68,8'd76,8'd20};
            mem_ROMWRAP[549] = {8'd69,8'd77,8'd20};
            mem_ROMWRAP[550] = {8'd70,8'd78,8'd20};
            mem_ROMWRAP[551] = {8'd71,8'd79,8'd20};
            mem_ROMWRAP[552] = {8'd80,8'd88,8'd21};
            mem_ROMWRAP[553] = {8'd81,8'd89,8'd21};
            mem_ROMWRAP[554] = {8'd82,8'd90,8'd21};
            mem_ROMWRAP[555] = {8'd83,8'd91,8'd21};
            mem_ROMWRAP[556] = {8'd84,8'd92,8'd21};
            mem_ROMWRAP[557] = {8'd85,8'd93,8'd21};
            mem_ROMWRAP[558] = {8'd86,8'd94,8'd21};
            mem_ROMWRAP[559] = {8'd87,8'd95,8'd21};
            mem_ROMWRAP[560] = {8'd96,8'd104,8'd22};
            mem_ROMWRAP[561] = {8'd97,8'd105,8'd22};
            mem_ROMWRAP[562] = {8'd98,8'd106,8'd22};
            mem_ROMWRAP[563] = {8'd99,8'd107,8'd22};
            mem_ROMWRAP[564] = {8'd100,8'd108,8'd22};
            mem_ROMWRAP[565] = {8'd101,8'd109,8'd22};
            mem_ROMWRAP[566] = {8'd102,8'd110,8'd22};
            mem_ROMWRAP[567] = {8'd103,8'd111,8'd22};
            mem_ROMWRAP[568] = {8'd112,8'd120,8'd23};
            mem_ROMWRAP[569] = {8'd113,8'd121,8'd23};
            mem_ROMWRAP[570] = {8'd114,8'd122,8'd23};
            mem_ROMWRAP[571] = {8'd115,8'd123,8'd23};
            mem_ROMWRAP[572] = {8'd116,8'd124,8'd23};
            mem_ROMWRAP[573] = {8'd117,8'd125,8'd23};
            mem_ROMWRAP[574] = {8'd118,8'd126,8'd23};
            mem_ROMWRAP[575] = {8'd119,8'd127,8'd23};
            mem_ROMWRAP[576] = {8'd128,8'd136,8'd24};
            mem_ROMWRAP[577] = {8'd129,8'd137,8'd24};
            mem_ROMWRAP[578] = {8'd130,8'd138,8'd24};
            mem_ROMWRAP[579] = {8'd131,8'd139,8'd24};
            mem_ROMWRAP[580] = {8'd132,8'd140,8'd24};
            mem_ROMWRAP[581] = {8'd133,8'd141,8'd24};
            mem_ROMWRAP[582] = {8'd134,8'd142,8'd24};
            mem_ROMWRAP[583] = {8'd135,8'd143,8'd24};
            mem_ROMWRAP[584] = {8'd144,8'd152,8'd25};
            mem_ROMWRAP[585] = {8'd145,8'd153,8'd25};
            mem_ROMWRAP[586] = {8'd146,8'd154,8'd25};
            mem_ROMWRAP[587] = {8'd147,8'd155,8'd25};
            mem_ROMWRAP[588] = {8'd148,8'd156,8'd25};
            mem_ROMWRAP[589] = {8'd149,8'd157,8'd25};
            mem_ROMWRAP[590] = {8'd150,8'd158,8'd25};
            mem_ROMWRAP[591] = {8'd151,8'd159,8'd25};
            mem_ROMWRAP[592] = {8'd160,8'd168,8'd26};
            mem_ROMWRAP[593] = {8'd161,8'd169,8'd26};
            mem_ROMWRAP[594] = {8'd162,8'd170,8'd26};
            mem_ROMWRAP[595] = {8'd163,8'd171,8'd26};
            mem_ROMWRAP[596] = {8'd164,8'd172,8'd26};
            mem_ROMWRAP[597] = {8'd165,8'd173,8'd26};
            mem_ROMWRAP[598] = {8'd166,8'd174,8'd26};
            mem_ROMWRAP[599] = {8'd167,8'd175,8'd26};
            mem_ROMWRAP[600] = {8'd176,8'd184,8'd27};
            mem_ROMWRAP[601] = {8'd177,8'd185,8'd27};
            mem_ROMWRAP[602] = {8'd178,8'd186,8'd27};
            mem_ROMWRAP[603] = {8'd179,8'd187,8'd27};
            mem_ROMWRAP[604] = {8'd180,8'd188,8'd27};
            mem_ROMWRAP[605] = {8'd181,8'd189,8'd27};
            mem_ROMWRAP[606] = {8'd182,8'd190,8'd27};
            mem_ROMWRAP[607] = {8'd183,8'd191,8'd27};
            mem_ROMWRAP[608] = {8'd192,8'd200,8'd28};
            mem_ROMWRAP[609] = {8'd193,8'd201,8'd28};
            mem_ROMWRAP[610] = {8'd194,8'd202,8'd28};
            mem_ROMWRAP[611] = {8'd195,8'd203,8'd28};
            mem_ROMWRAP[612] = {8'd196,8'd204,8'd28};
            mem_ROMWRAP[613] = {8'd197,8'd205,8'd28};
            mem_ROMWRAP[614] = {8'd198,8'd206,8'd28};
            mem_ROMWRAP[615] = {8'd199,8'd207,8'd28};
            mem_ROMWRAP[616] = {8'd208,8'd216,8'd29};
            mem_ROMWRAP[617] = {8'd209,8'd217,8'd29};
            mem_ROMWRAP[618] = {8'd210,8'd218,8'd29};
            mem_ROMWRAP[619] = {8'd211,8'd219,8'd29};
            mem_ROMWRAP[620] = {8'd212,8'd220,8'd29};
            mem_ROMWRAP[621] = {8'd213,8'd221,8'd29};
            mem_ROMWRAP[622] = {8'd214,8'd222,8'd29};
            mem_ROMWRAP[623] = {8'd215,8'd223,8'd29};
            mem_ROMWRAP[624] = {8'd224,8'd232,8'd30};
            mem_ROMWRAP[625] = {8'd225,8'd233,8'd30};
            mem_ROMWRAP[626] = {8'd226,8'd234,8'd30};
            mem_ROMWRAP[627] = {8'd227,8'd235,8'd30};
            mem_ROMWRAP[628] = {8'd228,8'd236,8'd30};
            mem_ROMWRAP[629] = {8'd229,8'd237,8'd30};
            mem_ROMWRAP[630] = {8'd230,8'd238,8'd30};
            mem_ROMWRAP[631] = {8'd231,8'd239,8'd30};
            mem_ROMWRAP[632] = {8'd240,8'd248,8'd31};
            mem_ROMWRAP[633] = {8'd241,8'd249,8'd31};
            mem_ROMWRAP[634] = {8'd242,8'd250,8'd31};
            mem_ROMWRAP[635] = {8'd243,8'd251,8'd31};
            mem_ROMWRAP[636] = {8'd244,8'd252,8'd31};
            mem_ROMWRAP[637] = {8'd245,8'd253,8'd31};
            mem_ROMWRAP[638] = {8'd246,8'd254,8'd31};
            mem_ROMWRAP[639] = {8'd247,8'd255,8'd31};
            mem_ROMWRAP[640] = {8'd0,8'd4,8'd32};
            mem_ROMWRAP[641] = {8'd1,8'd5,8'd32};
            mem_ROMWRAP[642] = {8'd2,8'd6,8'd32};
            mem_ROMWRAP[643] = {8'd3,8'd7,8'd32};
            mem_ROMWRAP[644] = {8'd8,8'd12,8'd33};
            mem_ROMWRAP[645] = {8'd9,8'd13,8'd33};
            mem_ROMWRAP[646] = {8'd10,8'd14,8'd33};
            mem_ROMWRAP[647] = {8'd11,8'd15,8'd33};
            mem_ROMWRAP[648] = {8'd16,8'd20,8'd34};
            mem_ROMWRAP[649] = {8'd17,8'd21,8'd34};
            mem_ROMWRAP[650] = {8'd18,8'd22,8'd34};
            mem_ROMWRAP[651] = {8'd19,8'd23,8'd34};
            mem_ROMWRAP[652] = {8'd24,8'd28,8'd35};
            mem_ROMWRAP[653] = {8'd25,8'd29,8'd35};
            mem_ROMWRAP[654] = {8'd26,8'd30,8'd35};
            mem_ROMWRAP[655] = {8'd27,8'd31,8'd35};
            mem_ROMWRAP[656] = {8'd32,8'd36,8'd36};
            mem_ROMWRAP[657] = {8'd33,8'd37,8'd36};
            mem_ROMWRAP[658] = {8'd34,8'd38,8'd36};
            mem_ROMWRAP[659] = {8'd35,8'd39,8'd36};
            mem_ROMWRAP[660] = {8'd40,8'd44,8'd37};
            mem_ROMWRAP[661] = {8'd41,8'd45,8'd37};
            mem_ROMWRAP[662] = {8'd42,8'd46,8'd37};
            mem_ROMWRAP[663] = {8'd43,8'd47,8'd37};
            mem_ROMWRAP[664] = {8'd48,8'd52,8'd38};
            mem_ROMWRAP[665] = {8'd49,8'd53,8'd38};
            mem_ROMWRAP[666] = {8'd50,8'd54,8'd38};
            mem_ROMWRAP[667] = {8'd51,8'd55,8'd38};
            mem_ROMWRAP[668] = {8'd56,8'd60,8'd39};
            mem_ROMWRAP[669] = {8'd57,8'd61,8'd39};
            mem_ROMWRAP[670] = {8'd58,8'd62,8'd39};
            mem_ROMWRAP[671] = {8'd59,8'd63,8'd39};
            mem_ROMWRAP[672] = {8'd64,8'd68,8'd40};
            mem_ROMWRAP[673] = {8'd65,8'd69,8'd40};
            mem_ROMWRAP[674] = {8'd66,8'd70,8'd40};
            mem_ROMWRAP[675] = {8'd67,8'd71,8'd40};
            mem_ROMWRAP[676] = {8'd72,8'd76,8'd41};
            mem_ROMWRAP[677] = {8'd73,8'd77,8'd41};
            mem_ROMWRAP[678] = {8'd74,8'd78,8'd41};
            mem_ROMWRAP[679] = {8'd75,8'd79,8'd41};
            mem_ROMWRAP[680] = {8'd80,8'd84,8'd42};
            mem_ROMWRAP[681] = {8'd81,8'd85,8'd42};
            mem_ROMWRAP[682] = {8'd82,8'd86,8'd42};
            mem_ROMWRAP[683] = {8'd83,8'd87,8'd42};
            mem_ROMWRAP[684] = {8'd88,8'd92,8'd43};
            mem_ROMWRAP[685] = {8'd89,8'd93,8'd43};
            mem_ROMWRAP[686] = {8'd90,8'd94,8'd43};
            mem_ROMWRAP[687] = {8'd91,8'd95,8'd43};
            mem_ROMWRAP[688] = {8'd96,8'd100,8'd44};
            mem_ROMWRAP[689] = {8'd97,8'd101,8'd44};
            mem_ROMWRAP[690] = {8'd98,8'd102,8'd44};
            mem_ROMWRAP[691] = {8'd99,8'd103,8'd44};
            mem_ROMWRAP[692] = {8'd104,8'd108,8'd45};
            mem_ROMWRAP[693] = {8'd105,8'd109,8'd45};
            mem_ROMWRAP[694] = {8'd106,8'd110,8'd45};
            mem_ROMWRAP[695] = {8'd107,8'd111,8'd45};
            mem_ROMWRAP[696] = {8'd112,8'd116,8'd46};
            mem_ROMWRAP[697] = {8'd113,8'd117,8'd46};
            mem_ROMWRAP[698] = {8'd114,8'd118,8'd46};
            mem_ROMWRAP[699] = {8'd115,8'd119,8'd46};
            mem_ROMWRAP[700] = {8'd120,8'd124,8'd47};
            mem_ROMWRAP[701] = {8'd121,8'd125,8'd47};
            mem_ROMWRAP[702] = {8'd122,8'd126,8'd47};
            mem_ROMWRAP[703] = {8'd123,8'd127,8'd47};
            mem_ROMWRAP[704] = {8'd128,8'd132,8'd48};
            mem_ROMWRAP[705] = {8'd129,8'd133,8'd48};
            mem_ROMWRAP[706] = {8'd130,8'd134,8'd48};
            mem_ROMWRAP[707] = {8'd131,8'd135,8'd48};
            mem_ROMWRAP[708] = {8'd136,8'd140,8'd49};
            mem_ROMWRAP[709] = {8'd137,8'd141,8'd49};
            mem_ROMWRAP[710] = {8'd138,8'd142,8'd49};
            mem_ROMWRAP[711] = {8'd139,8'd143,8'd49};
            mem_ROMWRAP[712] = {8'd144,8'd148,8'd50};
            mem_ROMWRAP[713] = {8'd145,8'd149,8'd50};
            mem_ROMWRAP[714] = {8'd146,8'd150,8'd50};
            mem_ROMWRAP[715] = {8'd147,8'd151,8'd50};
            mem_ROMWRAP[716] = {8'd152,8'd156,8'd51};
            mem_ROMWRAP[717] = {8'd153,8'd157,8'd51};
            mem_ROMWRAP[718] = {8'd154,8'd158,8'd51};
            mem_ROMWRAP[719] = {8'd155,8'd159,8'd51};
            mem_ROMWRAP[720] = {8'd160,8'd164,8'd52};
            mem_ROMWRAP[721] = {8'd161,8'd165,8'd52};
            mem_ROMWRAP[722] = {8'd162,8'd166,8'd52};
            mem_ROMWRAP[723] = {8'd163,8'd167,8'd52};
            mem_ROMWRAP[724] = {8'd168,8'd172,8'd53};
            mem_ROMWRAP[725] = {8'd169,8'd173,8'd53};
            mem_ROMWRAP[726] = {8'd170,8'd174,8'd53};
            mem_ROMWRAP[727] = {8'd171,8'd175,8'd53};
            mem_ROMWRAP[728] = {8'd176,8'd180,8'd54};
            mem_ROMWRAP[729] = {8'd177,8'd181,8'd54};
            mem_ROMWRAP[730] = {8'd178,8'd182,8'd54};
            mem_ROMWRAP[731] = {8'd179,8'd183,8'd54};
            mem_ROMWRAP[732] = {8'd184,8'd188,8'd55};
            mem_ROMWRAP[733] = {8'd185,8'd189,8'd55};
            mem_ROMWRAP[734] = {8'd186,8'd190,8'd55};
            mem_ROMWRAP[735] = {8'd187,8'd191,8'd55};
            mem_ROMWRAP[736] = {8'd192,8'd196,8'd56};
            mem_ROMWRAP[737] = {8'd193,8'd197,8'd56};
            mem_ROMWRAP[738] = {8'd194,8'd198,8'd56};
            mem_ROMWRAP[739] = {8'd195,8'd199,8'd56};
            mem_ROMWRAP[740] = {8'd200,8'd204,8'd57};
            mem_ROMWRAP[741] = {8'd201,8'd205,8'd57};
            mem_ROMWRAP[742] = {8'd202,8'd206,8'd57};
            mem_ROMWRAP[743] = {8'd203,8'd207,8'd57};
            mem_ROMWRAP[744] = {8'd208,8'd212,8'd58};
            mem_ROMWRAP[745] = {8'd209,8'd213,8'd58};
            mem_ROMWRAP[746] = {8'd210,8'd214,8'd58};
            mem_ROMWRAP[747] = {8'd211,8'd215,8'd58};
            mem_ROMWRAP[748] = {8'd216,8'd220,8'd59};
            mem_ROMWRAP[749] = {8'd217,8'd221,8'd59};
            mem_ROMWRAP[750] = {8'd218,8'd222,8'd59};
            mem_ROMWRAP[751] = {8'd219,8'd223,8'd59};
            mem_ROMWRAP[752] = {8'd224,8'd228,8'd60};
            mem_ROMWRAP[753] = {8'd225,8'd229,8'd60};
            mem_ROMWRAP[754] = {8'd226,8'd230,8'd60};
            mem_ROMWRAP[755] = {8'd227,8'd231,8'd60};
            mem_ROMWRAP[756] = {8'd232,8'd236,8'd61};
            mem_ROMWRAP[757] = {8'd233,8'd237,8'd61};
            mem_ROMWRAP[758] = {8'd234,8'd238,8'd61};
            mem_ROMWRAP[759] = {8'd235,8'd239,8'd61};
            mem_ROMWRAP[760] = {8'd240,8'd244,8'd62};
            mem_ROMWRAP[761] = {8'd241,8'd245,8'd62};
            mem_ROMWRAP[762] = {8'd242,8'd246,8'd62};
            mem_ROMWRAP[763] = {8'd243,8'd247,8'd62};
            mem_ROMWRAP[764] = {8'd248,8'd252,8'd63};
            mem_ROMWRAP[765] = {8'd249,8'd253,8'd63};
            mem_ROMWRAP[766] = {8'd250,8'd254,8'd63};
            mem_ROMWRAP[767] = {8'd251,8'd255,8'd63};
            mem_ROMWRAP[768] = {8'd0,8'd2,8'd64};
            mem_ROMWRAP[769] = {8'd1,8'd3,8'd64};
            mem_ROMWRAP[770] = {8'd4,8'd6,8'd65};
            mem_ROMWRAP[771] = {8'd5,8'd7,8'd65};
            mem_ROMWRAP[772] = {8'd8,8'd10,8'd66};
            mem_ROMWRAP[773] = {8'd9,8'd11,8'd66};
            mem_ROMWRAP[774] = {8'd12,8'd14,8'd67};
            mem_ROMWRAP[775] = {8'd13,8'd15,8'd67};
            mem_ROMWRAP[776] = {8'd16,8'd18,8'd68};
            mem_ROMWRAP[777] = {8'd17,8'd19,8'd68};
            mem_ROMWRAP[778] = {8'd20,8'd22,8'd69};
            mem_ROMWRAP[779] = {8'd21,8'd23,8'd69};
            mem_ROMWRAP[780] = {8'd24,8'd26,8'd70};
            mem_ROMWRAP[781] = {8'd25,8'd27,8'd70};
            mem_ROMWRAP[782] = {8'd28,8'd30,8'd71};
            mem_ROMWRAP[783] = {8'd29,8'd31,8'd71};
            mem_ROMWRAP[784] = {8'd32,8'd34,8'd72};
            mem_ROMWRAP[785] = {8'd33,8'd35,8'd72};
            mem_ROMWRAP[786] = {8'd36,8'd38,8'd73};
            mem_ROMWRAP[787] = {8'd37,8'd39,8'd73};
            mem_ROMWRAP[788] = {8'd40,8'd42,8'd74};
            mem_ROMWRAP[789] = {8'd41,8'd43,8'd74};
            mem_ROMWRAP[790] = {8'd44,8'd46,8'd75};
            mem_ROMWRAP[791] = {8'd45,8'd47,8'd76};
            mem_ROMWRAP[792] = {8'd48,8'd50,8'd76};
            mem_ROMWRAP[793] = {8'd49,8'd51,8'd76};
            mem_ROMWRAP[794] = {8'd52,8'd54,8'd77};
            mem_ROMWRAP[795] = {8'd53,8'd55,8'd77};
            mem_ROMWRAP[796] = {8'd56,8'd58,8'd78};
            mem_ROMWRAP[797] = {8'd57,8'd59,8'd78};
            mem_ROMWRAP[798] = {8'd60,8'd62,8'd79};
            mem_ROMWRAP[799] = {8'd61,8'd63,8'd79};
            mem_ROMWRAP[800] = {8'd64,8'd66,8'd80};
            mem_ROMWRAP[801] = {8'd65,8'd67,8'd80};
            mem_ROMWRAP[802] = {8'd68,8'd70,8'd81};
            mem_ROMWRAP[803] = {8'd69,8'd71,8'd81};
            mem_ROMWRAP[804] = {8'd72,8'd74,8'd82};
            mem_ROMWRAP[805] = {8'd73,8'd75,8'd82};
            mem_ROMWRAP[806] = {8'd76,8'd78,8'd83};
            mem_ROMWRAP[807] = {8'd77,8'd79,8'd83};
            mem_ROMWRAP[808] = {8'd80,8'd82,8'd84};
            mem_ROMWRAP[809] = {8'd81,8'd83,8'd84};
            mem_ROMWRAP[810] = {8'd84,8'd86,8'd85};
            mem_ROMWRAP[811] = {8'd85,8'd87,8'd85};
            mem_ROMWRAP[812] = {8'd88,8'd90,8'd86};
            mem_ROMWRAP[813] = {8'd89,8'd91,8'd86};
            mem_ROMWRAP[814] = {8'd92,8'd94,8'd87};
            mem_ROMWRAP[815] = {8'd93,8'd95,8'd87};
            mem_ROMWRAP[816] = {8'd96,8'd98,8'd88};
            mem_ROMWRAP[817] = {8'd97,8'd99,8'd88};
            mem_ROMWRAP[818] = {8'd100,8'd102,8'd89};
            mem_ROMWRAP[819] = {8'd101,8'd103,8'd89};
            mem_ROMWRAP[820] = {8'd104,8'd106,8'd90};
            mem_ROMWRAP[821] = {8'd105,8'd107,8'd90};
            mem_ROMWRAP[822] = {8'd108,8'd110,8'd91};
            mem_ROMWRAP[823] = {8'd109,8'd111,8'd91};
            mem_ROMWRAP[824] = {8'd112,8'd114,8'd92};
            mem_ROMWRAP[825] = {8'd113,8'd115,8'd92};
            mem_ROMWRAP[826] = {8'd116,8'd118,8'd93};
            mem_ROMWRAP[827] = {8'd117,8'd119,8'd93};
            mem_ROMWRAP[828] = {8'd120,8'd122,8'd94};
            mem_ROMWRAP[829] = {8'd121,8'd123,8'd94};
            mem_ROMWRAP[830] = {8'd124,8'd126,8'd95};
            mem_ROMWRAP[831] = {8'd125,8'd127,8'd95};
            mem_ROMWRAP[832] = {8'd128,8'd130,8'd96};
            mem_ROMWRAP[833] = {8'd129,8'd131,8'd96};
            mem_ROMWRAP[834] = {8'd132,8'd134,8'd97};
            mem_ROMWRAP[835] = {8'd133,8'd135,8'd97};
            mem_ROMWRAP[836] = {8'd136,8'd138,8'd98};
            mem_ROMWRAP[837] = {8'd137,8'd139,8'd98};
            mem_ROMWRAP[838] = {8'd140,8'd142,8'd99};
            mem_ROMWRAP[839] = {8'd141,8'd143,8'd99};
            mem_ROMWRAP[840] = {8'd144,8'd146,8'd100};
            mem_ROMWRAP[841] = {8'd145,8'd147,8'd100};
            mem_ROMWRAP[842] = {8'd148,8'd150,8'd101};
            mem_ROMWRAP[843] = {8'd149,8'd151,8'd101};
            mem_ROMWRAP[844] = {8'd152,8'd154,8'd102};
            mem_ROMWRAP[845] = {8'd153,8'd155,8'd102};
            mem_ROMWRAP[846] = {8'd156,8'd158,8'd103};
            mem_ROMWRAP[847] = {8'd157,8'd159,8'd103};
            mem_ROMWRAP[848] = {8'd160,8'd162,8'd104};
            mem_ROMWRAP[849] = {8'd161,8'd163,8'd104};
            mem_ROMWRAP[850] = {8'd164,8'd166,8'd105};
            mem_ROMWRAP[851] = {8'd165,8'd167,8'd105};
            mem_ROMWRAP[852] = {8'd168,8'd170,8'd106};
            mem_ROMWRAP[853] = {8'd169,8'd171,8'd106};
            mem_ROMWRAP[854] = {8'd172,8'd174,8'd107};
            mem_ROMWRAP[855] = {8'd173,8'd175,8'd107};
            mem_ROMWRAP[856] = {8'd176,8'd178,8'd108};
            mem_ROMWRAP[857] = {8'd177,8'd179,8'd108};
            mem_ROMWRAP[858] = {8'd180,8'd182,8'd109};
            mem_ROMWRAP[859] = {8'd181,8'd183,8'd109};
            mem_ROMWRAP[860] = {8'd184,8'd186,8'd110};
            mem_ROMWRAP[861] = {8'd185,8'd187,8'd110};
            mem_ROMWRAP[862] = {8'd188,8'd190,8'd111};
            mem_ROMWRAP[863] = {8'd189,8'd191,8'd111};
            mem_ROMWRAP[864] = {8'd192,8'd194,8'd112};
            mem_ROMWRAP[865] = {8'd193,8'd195,8'd112};
            mem_ROMWRAP[866] = {8'd196,8'd198,8'd113};
            mem_ROMWRAP[867] = {8'd197,8'd199,8'd113};
            mem_ROMWRAP[868] = {8'd200,8'd202,8'd114};
            mem_ROMWRAP[869] = {8'd201,8'd203,8'd114};
            mem_ROMWRAP[870] = {8'd204,8'd206,8'd115};
            mem_ROMWRAP[871] = {8'd205,8'd207,8'd115};
            mem_ROMWRAP[872] = {8'd208,8'd210,8'd116};
            mem_ROMWRAP[873] = {8'd209,8'd211,8'd116};
            mem_ROMWRAP[874] = {8'd212,8'd214,8'd117};
            mem_ROMWRAP[875] = {8'd213,8'd215,8'd117};
            mem_ROMWRAP[876] = {8'd216,8'd218,8'd118};
            mem_ROMWRAP[877] = {8'd217,8'd219,8'd118};
            mem_ROMWRAP[878] = {8'd220,8'd222,8'd119};
            mem_ROMWRAP[879] = {8'd221,8'd223,8'd119};
            mem_ROMWRAP[880] = {8'd224,8'd226,8'd120};
            mem_ROMWRAP[881] = {8'd225,8'd227,8'd120};
            mem_ROMWRAP[882] = {8'd228,8'd230,8'd121};
            mem_ROMWRAP[883] = {8'd229,8'd231,8'd121};
            mem_ROMWRAP[884] = {8'd232,8'd234,8'd122};
            mem_ROMWRAP[885] = {8'd233,8'd235,8'd122};
            mem_ROMWRAP[886] = {8'd236,8'd238,8'd123};
            mem_ROMWRAP[887] = {8'd237,8'd239,8'd123};
            mem_ROMWRAP[888] = {8'd240,8'd242,8'd124};
            mem_ROMWRAP[889] = {8'd241,8'd243,8'd124};
            mem_ROMWRAP[890] = {8'd244,8'd246,8'd125};
            mem_ROMWRAP[891] = {8'd245,8'd247,8'd125};
            mem_ROMWRAP[892] = {8'd248,8'd250,8'd126};
            mem_ROMWRAP[893] = {8'd249,8'd251,8'd126};
            mem_ROMWRAP[894] = {8'd252,8'd254,8'd127};
            mem_ROMWRAP[895] = {8'd253,8'd255,8'd127};
	end

	always @(posedge clk)
	begin
		a <= mem_ROMWRAP[address1];
	end  
endmodule

