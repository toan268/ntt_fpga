
module soc_system (
	button_pio_external_connection_export,
	clk_clk,
	dipsw_pio_external_connection_export,
	hps_0_f2h_cold_reset_req_reset_n,
	hps_0_f2h_debug_reset_req_reset_n,
	hps_0_f2h_stm_hw_events_stm_hwevents,
	hps_0_f2h_warm_reset_req_reset_n,
	hps_0_h2f_reset_reset_n,
	hps_0_hps_io_hps_io_emac1_inst_TX_CLK,
	hps_0_hps_io_hps_io_emac1_inst_TXD0,
	hps_0_hps_io_hps_io_emac1_inst_TXD1,
	hps_0_hps_io_hps_io_emac1_inst_TXD2,
	hps_0_hps_io_hps_io_emac1_inst_TXD3,
	hps_0_hps_io_hps_io_emac1_inst_RXD0,
	hps_0_hps_io_hps_io_emac1_inst_MDIO,
	hps_0_hps_io_hps_io_emac1_inst_MDC,
	hps_0_hps_io_hps_io_emac1_inst_RX_CTL,
	hps_0_hps_io_hps_io_emac1_inst_TX_CTL,
	hps_0_hps_io_hps_io_emac1_inst_RX_CLK,
	hps_0_hps_io_hps_io_emac1_inst_RXD1,
	hps_0_hps_io_hps_io_emac1_inst_RXD2,
	hps_0_hps_io_hps_io_emac1_inst_RXD3,
	hps_0_hps_io_hps_io_qspi_inst_IO0,
	hps_0_hps_io_hps_io_qspi_inst_IO1,
	hps_0_hps_io_hps_io_qspi_inst_IO2,
	hps_0_hps_io_hps_io_qspi_inst_IO3,
	hps_0_hps_io_hps_io_qspi_inst_SS0,
	hps_0_hps_io_hps_io_qspi_inst_CLK,
	hps_0_hps_io_hps_io_sdio_inst_CMD,
	hps_0_hps_io_hps_io_sdio_inst_D0,
	hps_0_hps_io_hps_io_sdio_inst_D1,
	hps_0_hps_io_hps_io_sdio_inst_CLK,
	hps_0_hps_io_hps_io_sdio_inst_D2,
	hps_0_hps_io_hps_io_sdio_inst_D3,
	hps_0_hps_io_hps_io_usb1_inst_D0,
	hps_0_hps_io_hps_io_usb1_inst_D1,
	hps_0_hps_io_hps_io_usb1_inst_D2,
	hps_0_hps_io_hps_io_usb1_inst_D3,
	hps_0_hps_io_hps_io_usb1_inst_D4,
	hps_0_hps_io_hps_io_usb1_inst_D5,
	hps_0_hps_io_hps_io_usb1_inst_D6,
	hps_0_hps_io_hps_io_usb1_inst_D7,
	hps_0_hps_io_hps_io_usb1_inst_CLK,
	hps_0_hps_io_hps_io_usb1_inst_STP,
	hps_0_hps_io_hps_io_usb1_inst_DIR,
	hps_0_hps_io_hps_io_usb1_inst_NXT,
	hps_0_hps_io_hps_io_spim0_inst_CLK,
	hps_0_hps_io_hps_io_spim0_inst_MOSI,
	hps_0_hps_io_hps_io_spim0_inst_MISO,
	hps_0_hps_io_hps_io_spim0_inst_SS0,
	hps_0_hps_io_hps_io_spim1_inst_CLK,
	hps_0_hps_io_hps_io_spim1_inst_MOSI,
	hps_0_hps_io_hps_io_spim1_inst_MISO,
	hps_0_hps_io_hps_io_spim1_inst_SS0,
	hps_0_hps_io_hps_io_uart0_inst_RX,
	hps_0_hps_io_hps_io_uart0_inst_TX,
	hps_0_hps_io_hps_io_i2c0_inst_SDA,
	hps_0_hps_io_hps_io_i2c0_inst_SCL,
	hps_0_hps_io_hps_io_i2c1_inst_SDA,
	hps_0_hps_io_hps_io_i2c1_inst_SCL,
	hps_0_hps_io_hps_io_gpio_inst_GPIO09,
	hps_0_hps_io_hps_io_gpio_inst_GPIO35,
	hps_0_hps_io_hps_io_gpio_inst_GPIO37,
	hps_0_hps_io_hps_io_gpio_inst_GPIO40,
	hps_0_hps_io_hps_io_gpio_inst_GPIO41,
	hps_0_hps_io_hps_io_gpio_inst_GPIO44,
	hps_0_hps_io_hps_io_gpio_inst_GPIO48,
	hps_0_hps_io_hps_io_gpio_inst_GPIO53,
	hps_0_hps_io_hps_io_gpio_inst_GPIO54,
	hps_0_hps_io_hps_io_gpio_inst_GPIO61,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	reset_reset_n,
	f2h_sdram0_data_address,
	f2h_sdram0_data_read,
	f2h_sdram0_data_readdata,
	f2h_sdram0_data_write,
	f2h_sdram0_data_writedata,
	f2h_sdram0_data_readdatavalid,
	f2h_sdram0_data_waitrequest,
	f2h_sdram0_data_byteenable,
	f2h_sdram0_data_burstcount,
	f2h_sdram0_cntl_read,
	f2h_sdram0_cntl_readdata,
	f2h_sdram0_cntl_write,
	f2h_sdram0_cntl_writedata,
	f2h_sdram0_cntl_byteenable,
	slave_template_0_user_interface_dataout_0,
	slave_template_0_user_interface_dataout_1,
	slave_template_0_user_interface_dataout_2,
	slave_template_0_user_interface_dataout_3,
	slave_template_0_user_interface_dataout_4,
	slave_template_0_user_interface_dataout_5,
	slave_template_0_user_interface_dataout_6,
	slave_template_0_user_interface_dataout_7,
	slave_template_0_user_interface_dataout_8,
	slave_template_0_user_interface_dataout_9,
	slave_template_0_user_interface_dataout_10,
	slave_template_0_user_interface_dataout_11,
	slave_template_0_user_interface_dataout_12,
	slave_template_0_user_interface_dataout_13,
	slave_template_0_user_interface_dataout_14,
	slave_template_0_user_interface_dataout_15,
	slave_template_0_user_interface_datain_0,
	slave_template_0_user_interface_datain_1,
	slave_template_0_user_interface_datain_2,
	slave_template_0_user_interface_datain_3,
	slave_template_0_user_interface_datain_4,
	slave_template_0_user_interface_datain_5,
	slave_template_0_user_interface_datain_6,
	slave_template_0_user_interface_datain_7,
	slave_template_0_user_interface_datain_8,
	slave_template_0_user_interface_datain_9,
	slave_template_0_user_interface_datain_10,
	slave_template_0_user_interface_datain_11,
	slave_template_0_user_interface_datain_12,
	slave_template_0_user_interface_datain_13,
	slave_template_0_user_interface_datain_14,
	slave_template_0_user_interface_datain_15);	

	input	[3:0]	button_pio_external_connection_export;
	input		clk_clk;
	input	[9:0]	dipsw_pio_external_connection_export;
	input		hps_0_f2h_cold_reset_req_reset_n;
	input		hps_0_f2h_debug_reset_req_reset_n;
	input	[27:0]	hps_0_f2h_stm_hw_events_stm_hwevents;
	input		hps_0_f2h_warm_reset_req_reset_n;
	output		hps_0_h2f_reset_reset_n;
	output		hps_0_hps_io_hps_io_emac1_inst_TX_CLK;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD0;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD1;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD2;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD3;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD0;
	inout		hps_0_hps_io_hps_io_emac1_inst_MDIO;
	output		hps_0_hps_io_hps_io_emac1_inst_MDC;
	input		hps_0_hps_io_hps_io_emac1_inst_RX_CTL;
	output		hps_0_hps_io_hps_io_emac1_inst_TX_CTL;
	input		hps_0_hps_io_hps_io_emac1_inst_RX_CLK;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD1;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD2;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD3;
	inout		hps_0_hps_io_hps_io_qspi_inst_IO0;
	inout		hps_0_hps_io_hps_io_qspi_inst_IO1;
	inout		hps_0_hps_io_hps_io_qspi_inst_IO2;
	inout		hps_0_hps_io_hps_io_qspi_inst_IO3;
	output		hps_0_hps_io_hps_io_qspi_inst_SS0;
	output		hps_0_hps_io_hps_io_qspi_inst_CLK;
	inout		hps_0_hps_io_hps_io_sdio_inst_CMD;
	inout		hps_0_hps_io_hps_io_sdio_inst_D0;
	inout		hps_0_hps_io_hps_io_sdio_inst_D1;
	output		hps_0_hps_io_hps_io_sdio_inst_CLK;
	inout		hps_0_hps_io_hps_io_sdio_inst_D2;
	inout		hps_0_hps_io_hps_io_sdio_inst_D3;
	inout		hps_0_hps_io_hps_io_usb1_inst_D0;
	inout		hps_0_hps_io_hps_io_usb1_inst_D1;
	inout		hps_0_hps_io_hps_io_usb1_inst_D2;
	inout		hps_0_hps_io_hps_io_usb1_inst_D3;
	inout		hps_0_hps_io_hps_io_usb1_inst_D4;
	inout		hps_0_hps_io_hps_io_usb1_inst_D5;
	inout		hps_0_hps_io_hps_io_usb1_inst_D6;
	inout		hps_0_hps_io_hps_io_usb1_inst_D7;
	input		hps_0_hps_io_hps_io_usb1_inst_CLK;
	output		hps_0_hps_io_hps_io_usb1_inst_STP;
	input		hps_0_hps_io_hps_io_usb1_inst_DIR;
	input		hps_0_hps_io_hps_io_usb1_inst_NXT;
	output		hps_0_hps_io_hps_io_spim0_inst_CLK;
	output		hps_0_hps_io_hps_io_spim0_inst_MOSI;
	input		hps_0_hps_io_hps_io_spim0_inst_MISO;
	output		hps_0_hps_io_hps_io_spim0_inst_SS0;
	output		hps_0_hps_io_hps_io_spim1_inst_CLK;
	output		hps_0_hps_io_hps_io_spim1_inst_MOSI;
	input		hps_0_hps_io_hps_io_spim1_inst_MISO;
	output		hps_0_hps_io_hps_io_spim1_inst_SS0;
	input		hps_0_hps_io_hps_io_uart0_inst_RX;
	output		hps_0_hps_io_hps_io_uart0_inst_TX;
	inout		hps_0_hps_io_hps_io_i2c0_inst_SDA;
	inout		hps_0_hps_io_hps_io_i2c0_inst_SCL;
	inout		hps_0_hps_io_hps_io_i2c1_inst_SDA;
	inout		hps_0_hps_io_hps_io_i2c1_inst_SCL;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO09;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO35;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO37;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO40;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO41;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO44;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO48;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO53;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO54;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO61;
	output	[14:0]	memory_mem_a;
	output	[2:0]	memory_mem_ba;
	output		memory_mem_ck;
	output		memory_mem_ck_n;
	output		memory_mem_cke;
	output		memory_mem_cs_n;
	output		memory_mem_ras_n;
	output		memory_mem_cas_n;
	output		memory_mem_we_n;
	output		memory_mem_reset_n;
	inout	[31:0]	memory_mem_dq;
	inout	[3:0]	memory_mem_dqs;
	inout	[3:0]	memory_mem_dqs_n;
	output		memory_mem_odt;
	output	[3:0]	memory_mem_dm;
	input		memory_oct_rzqin;
	input		reset_reset_n;
	input	[25:0]	f2h_sdram0_data_address;
	input		f2h_sdram0_data_read;
	output	[63:0]	f2h_sdram0_data_readdata;
	input		f2h_sdram0_data_write;
	input	[63:0]	f2h_sdram0_data_writedata;
	output		f2h_sdram0_data_readdatavalid;
	output		f2h_sdram0_data_waitrequest;
	input	[7:0]	f2h_sdram0_data_byteenable;
	input	[0:0]	f2h_sdram0_data_burstcount;
	input		f2h_sdram0_cntl_read;
	output	[63:0]	f2h_sdram0_cntl_readdata;
	input		f2h_sdram0_cntl_write;
	input	[63:0]	f2h_sdram0_cntl_writedata;
	input	[7:0]	f2h_sdram0_cntl_byteenable;
	output	[31:0]	slave_template_0_user_interface_dataout_0;
	output	[31:0]	slave_template_0_user_interface_dataout_1;
	output	[31:0]	slave_template_0_user_interface_dataout_2;
	output	[31:0]	slave_template_0_user_interface_dataout_3;
	output	[31:0]	slave_template_0_user_interface_dataout_4;
	output	[31:0]	slave_template_0_user_interface_dataout_5;
	output	[31:0]	slave_template_0_user_interface_dataout_6;
	output	[31:0]	slave_template_0_user_interface_dataout_7;
	output	[31:0]	slave_template_0_user_interface_dataout_8;
	output	[31:0]	slave_template_0_user_interface_dataout_9;
	output	[31:0]	slave_template_0_user_interface_dataout_10;
	output	[31:0]	slave_template_0_user_interface_dataout_11;
	output	[31:0]	slave_template_0_user_interface_dataout_12;
	output	[31:0]	slave_template_0_user_interface_dataout_13;
	output	[31:0]	slave_template_0_user_interface_dataout_14;
	output	[31:0]	slave_template_0_user_interface_dataout_15;
	input	[31:0]	slave_template_0_user_interface_datain_0;
	input	[31:0]	slave_template_0_user_interface_datain_1;
	input	[31:0]	slave_template_0_user_interface_datain_2;
	input	[31:0]	slave_template_0_user_interface_datain_3;
	input	[31:0]	slave_template_0_user_interface_datain_4;
	input	[31:0]	slave_template_0_user_interface_datain_5;
	input	[31:0]	slave_template_0_user_interface_datain_6;
	input	[31:0]	slave_template_0_user_interface_datain_7;
	input	[31:0]	slave_template_0_user_interface_datain_8;
	input	[31:0]	slave_template_0_user_interface_datain_9;
	input	[31:0]	slave_template_0_user_interface_datain_10;
	input	[31:0]	slave_template_0_user_interface_datain_11;
	input	[31:0]	slave_template_0_user_interface_datain_12;
	input	[31:0]	slave_template_0_user_interface_datain_13;
	input	[31:0]	slave_template_0_user_interface_datain_14;
	input	[31:0]	slave_template_0_user_interface_datain_15;
endmodule
